library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all ;

package IP_CORES is

  

end IP_CORES;
